Hanging branch
.circuit
V1 GND n1 dc 5
R1 GND n2 dc 5
R2 n2 n1 5
R4 n2 n3 5
V2 n3 n4 dc 10
.end