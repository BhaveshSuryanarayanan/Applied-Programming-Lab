Shorted Resistor 
.circuit
V1 n1 GND dc 5
R1 n1 n2 5
R2 GND n2 5
R3 n1 n1 5

.end